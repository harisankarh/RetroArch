BSV1        4  FCS�4  U&      ?  PC     [�A      P      %X       Y      �S      �RAM     dU � /�E �� t   i    �             �L     � �   ��q��� "        $  �' @�             P��   ��               ��        %                                                     	�  �����            � �  ****    � V���	������    � �                   ��  p0                   ��    �   � * "                                                              �������������������������������f�
{�� ������9�6Խ���ޮ��� ���[��
�b> T�
��
 
��
 �
��
�R�!�
��
 �
�rB�
��
��
 b< L�
 �
�
��
��
��
 R��
 �
��
�b>�
��
 �
�R�^�
��
��
 �
��
 �
�
 �
��
��
 b<�
 �
��
�R�V�
��
 �
�rB S�
��
�
 �
��
 �
�R�)�
��
��
 R�N�
 �
�                        dd                        U                                                                                                                                            _               �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             ! !+#"#* TT/'&'.TT       QQQQ   			
QQQ        ! +#"#"#TT/'&'&'        QQ;QQ  Q QQ QQ99                                UUU      U            ����                                    UU              P      �Z  ��           $  ����� 6:>_[[����'ë'˪'� '�P'�U'�P'��                                                                                                                                       )(0!076 &  �     ������������������������=   JAMM    IQLB       ICoa       ICou   ����TSBS   �6	    �	  NTAR          O     O  O   O   O        O O O   O O  O  O    O  O    O O O O   O O O     ��      ��       O   O   O  ������ ������  O   O          ������� �������    O           ����������������   O           ����� ������� ��       O                  �             454545454564545456454454    7898989:989:7898989:78987898    ;<===<=;=<=>;<===<=>;<==;<==    ^_2_22_22_^_^_2_2_^_^_2_^_2_            XYZ[XYZ[XYZ[XYZ[XYZ[XYZ[XYZ[    ����	
	
	
	
��������XYZ[XYZ[XYZ[��������	
	
	
	
	
	
	
����������������������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                �����������������       �PPPPPPP�UUUUPPP�����UUU��������               O O  O                    O O O    O  O                  O O O   O     ��                   O   O  ������                          ������                         �������                        ����� ��                                                5454545454545456                989:989:989:989:                =<=;=<=;=<=;=<=>                22_222_222_22_^_                                                XYZ[XYZ[XYZ[XYZ[                                	
	
 !!"	
                &01'                &01'                #$$%                	
	
                                XYZ[XYZ[                                ��������                ��������                ����������������                ����������������                                                                                ����    ����            PPPP    UU�U    PUUP    ����            PRAM    )(0!0 7 6  &   SPRA   
��
��
��
 R��
 �
��
�b>�
��
 �
�R�^�
��
��
 �
��
 �
�
 �
��
��
 b<�
 �
��
�R�V�
��
 �
�rB S�
��
�
 �
��
 �
�R�)�
��
��
 R�N�
 �
��
�b> T�
��
 
��
 �
��
�R�!�
��
 �
�rB�
��
��
 b< L�
 �
�PPUR   �@ KOOK   DEAD    PSPL    XOFF    VTOG    RADD   �TADD   �VBUF    PGEN   �   JYRB   JOYS       LSTS    �  FHCN   �[  FCNT    PSG    ����g	0ENCH   IQFM   NREG   ,ZTRIM    TRIC   E0SP   E1SP   E2SP    E0MO   E1MO   E2MO   E0D1   E1D1   E2D1   E0DV   E1DV   E2DV   LEN0   �   LEN1   �   LEN2   �   LEN3   �   SWEE     CRF1   �   CRF2   �   SWCT   SIRQ   �5ACC      5BIT   5ADD   Q|  5SIZ       5SHF    5VDM    5VSP    5SZL   5ADL   �5FMT   RWDA      CHRR     .24,۰ 1.,<�O ����B�������~�� 0 )>���g? 8!!!!>|�����> 0!9!c8|�����c !!!!�����o> ))!c�������c ?  >  ������� ?  >  ������� 8!!  g�������g�����[>�����><Z��ۥ[><fۥ��g>             " A     AAA"         88      ( 8       (            >:     .>&      >           <~~     <nNzf<     ~~<         <~��    <~����b<    ��~<        t�y    t<̅~��h    ���h    $V(
, <^4<8$8N $0<0V<
<8   ��[�z   �R��1    /    4b$<B��,^<<~��������~ ������~ 4b$����,^<����������� ������� 4b$����,^<����������� ������� 4b$����,^<����������� ������� 4b$����,^<����������� ������� 4b$����,^<����������� �������  5.N 69q��>�f3����y?�F���Z����KO�?���%��|�ے���  (;  /&~���o}{CC���PCg  ������  ������t��䨰p��~|xА , 3^]����g?ac�?	�y? � ����] ��� #����Zv�'?�o�������*Dy�6|I���X�!�(Ya��~�����$h��H$�<x���x<d��.#g�����`@@�    ����     �08���� ����|�v"		~>     	 8ĊB�����������L��p ��������F>     �z>                     ���     ���                           	      ?ww���� HH������@@3��?                     p�     p����xv���ތ��y~�L��00���������<       <       #!0�=>?���1}F� ��߻Ń ���o�������Ё�n/���p���ߋ�p    � @�    ����@ `�@�  ������  <r�����h<~�����wD_tf6{`Ky=          ?<1338?7><<?   =�o   3��������??a��#� |Ƃ:|�~ |��Ƃ��~X~�s�}9�������  ��   ����~F��>��<��^F���    s�    ��A�+_/���:Ԡ� �          	
6<6;0:  !���  ?��d�  �@  P� ��@            @ ��    @ ��  
0�     
0�                        :"e   >?{�gyw��]�񙏌 ���B<   ���~<                   �B����Ã����ġ<`� ������  ��@H�4 ���Ȝ,Ĥ8�    �|��    b��
  ~��   @@@@ @@ @@@@ @@                  |�r�  |�n�($�d$8<��� E��{��k�������__/    a`0                     s�s�F= n���=                 ��3��� �?���      8T      8l��<���������                ��x���E����  
/	  8	      $      <<?]W47w}�uߟ�sWW�����������@ ��b���� /__ 2c`]]'-bb:3� �����<���` p�윖�o�y�tzz����  ������  ��@@�` �X&	����z? 0L~�x� <|r�����ޯ'T������\o�
y���а��\�|t������ �܈H @�   �`�0Z�  ��Pj�9
  7       U�     U}��H     ˻H      
, 3^^]s=aacN# � ����x ���  ���������T4;?�??>                  ���@�  �*��p                                0(�I)"08��?>5F��D��~-�����~            �/_����ش���   <D|�?   <||�����*۴��;88�'O     ��     �R �|(�p����Ȑ`�  ?~�  6{�?  �z6   ~����   ~�~�����Á��~ <<�~�~   *  7"6???9 �h��� �����|������������9�   �����   �� 0��    �    8D����8|���}��_���A? ����>?~�������f��t�((p���@��  �����`��                 8x� (h�?O�=އ�_!? ��x?>? �@����� �����?����x��  �;���@��   ����   �EР�       �         %'&LH??;;:txHhp����xxxp����x����DD������||$$<<<<  :41  -;?~?OG!	"Y澞�>g���������������}y���   >?   !!=+2#7? "Y�^�� >g����\�<������t��r��  ��  `����~~9�_O/"Y�~>L�>g��������������������><|�����6<L�0 �������������??    #8    �������?``�       �       ������������<<<xx�<<,@H�a??6"��������``����p`����������@@�`����~����k�q�� �@����� ��������������    ����    �;�;�0      �0      1�"  � E	                             J1 /�1F	  "~n.�� >~r��tO5D�������    	=V   3yK%FUH�f|>�z\0`Q����6�_�9=���d�� � ��^�     0d        
�3    3	                                                 8D�r|r� 8|�~L~�                  _��  Z��        �������ݣ=�cx�    � А    ��0����B����x|����>� @��������� ��@������� �  ��@��  ���@  �����@                    �@���@  ������@@����� ���  ���                                                                                                                                                 �ϟ�??� �߿�� ?�����     �{. ������       � ������      � ������      
� .B!�   (H(4��A*��� KW��  LX��??�������t?�\,&33399��������^nv�������������{?1�3�?1�O���� ����� �3oG���<px�����ܮn����|<~�����������������          ��I�(c�	?[6; �M�Ų��Z�M8 �/ڛO��Q>�%$�  ���z��`@@  �@                    ��    ���X���� F�g�������7���������������ؤ������������xxx8���xxx8VL�����kn|�����l ������ ��????��Ga`��<��y���������~>���������`@OKKO�������� �  ��� �������  �������������OOKKP@������� ��� � ����� � �������������NNNNNNNN��������uuuuuuuu���������O�;w�<x� 0 ��9ܞ�����<  ��w�P����p0�����
�����`�c}����`X`�����?���?��~��c�c|����`P`��߇��?�?~�����������������?�?�?�?�����  �
۳��  � @    � �     ���   �f*�JU ��@�� �U�*D�  �TT        \       ;P@"	@*(J��4�1���110�jQ����""��$ydD�X DJJ ',%% %q`�Ed,Mip�`%Mi!5uuU@JPPP```BHPPP```�YF&Y&�&Y&d�R�����  �@@a" Q�d�&Q�� P�.IX�	�F�   
� �֊DHH QH(%%L	,V@
B� P�)J@�D��R(f�(�!Q�"�B��b�D$�2A�� � !�� @D	��0 @G��??�<�����d�����7399�������nd����������								��������Y&Y&Y&Y&Y&Y&Y&Y&                0�B��       x,�� $�$   �s�Ɠd�    `��I�L��     @	ɖ�VHɤ6�t!$       �CH+�       (�8�H�    @4 p'� 8�s �>�/v� ������  ��#G�  ��<x� �>��nw ���|~��5I�I�			ɤ6���$  ���@� ���v?�{l  �N�pi� ��@�  �<xp`R@������߿<������<�� @977��߿����>

�~���vz���0`@@P# �����ظ��66��~����6:� ����������� � ������?�����>xp`N3�����߿s����^�3o���E1�A�u�1���u�<r@C{���Ͽgo
|<������<��΀<aB;{���߿�yy�L����������uuuuu%�!�����%��3l;J��o;������ذ�� ���ؐ�� ?/MO� ������� �6�(pR����(pr�787-:���������8�h�������h�����"B ��ۻ��������B �����j���7s{<>� sqy<?�� ������ ������ NNNMBILP��������E5Z��" G7{��" ��x��� ������ {9;C`� y9����� ��\��   �����   ��uuu������Ac � ��ac � � � ���������� �  oO(���oo8���� � ����� � ����� ������ ����� ���� /;_O� ������� �0p�� �80��� � @;sw��߿�yqs>� ����>������RLIBAPLN���������80��X1A��7��{7G~.r���~������NNNNND[D�������߀ @0	���߳���>B�����>�������0`d@P/�����߿�(Pr*��pr*���JNT8@3����Իo'&
����������3�d&��'3�d&����̛&d�1��̛&d�37{8����9�x�����=�9��Ϝ;=���߼xs;	Ga� s?����� ��Zm��D ���o3�D u�u�E�5��u�ŵ5kks+�c� og?��� ���<|�  Ύ�<��  [@`TNNNN���������:�@� �;���� ޜ�x� ����� 18<� ������� ��hp�Ɔ ��xp�Ɔ �NGc� ������� ��<�� �<��� ;;�?�\ {{� ��,�� ������?���~�����������,�������
sf	 W�y�d<�0�` ;;�>�\ {z|� Col�?_/ ��/_/��JBA�����,0���0/0_�����[������h` ���@�`� �����   TZ4�    tu��1���    ����������      DJB���
@D@����
�$ �_�1��<�@@�������{�   � -�,�O����_(-TZ4�8?:0uu�og71����   �����
.�

Eeo�� ;;�?�\ c{{�π��    ߿��    � ��    ����    ??  ??     �f�j�`�`�f�o�`�`   ��    ���  �̚�2,� �ܺ�rl���������          <  ?            	    7c�Kǁ?����� ����`PP ����`PP `���� ��x|�p<    9   >( ??��p�|>_����������������  >���73  ��x8<<���ޔx\����ޔx\��p��  �����     ���   ����$2(0 trhhp   ���  ����  /0  ?0  264DI�???�
"+K����������������x<>  ������  ������      P��1!�Cs�������?O/�u7��������'	'	���[�v׾���������͏��_���������������Ѩ�����Ѩ   
#   
#?}럻i?}럻i����vҥ����vҥ����k�eX����k�eX    ���S�v׼����������+����������������o�������o�����������    �0�؟�� ��7`   ���?� ?�`�   ����o�  �~ �  `������ ��?   s��?����<0��@   ;g3O1O<<���$��@���$��@?  ?  @@@  �Y     �Y     tI�T0�@ tI�T0�@ �����n���������   O     0  ���  �������  ����  � �� �  ���   �0�؟�� ��7`   ���?� ?�`�   ����o�  �~ �  `������ ��?   s��?����<0��@   ��������        ���������   LATC   BUSC                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   